
--  _________  ________  ________        ________  _______   ________   _______   ________  ________  _________  ___  ________  ________           ________  _______   ________           ________  ________  ___  ___  ________                 ________  ___       _______   ________      
-- |\___   ___\\   __  \|\   __  \      |\   ____\|\  ___ \ |\   ___  \|\  ___ \ |\   __  \|\   __  \|\___   ___\\  \|\   __  \|\   ___  \        |\   ___ \|\  ___ \ |\   ____\         |\   ____\|\   __  \|\  \|\  \|\   ____\               |\   ____\|\  \     |\  ___ \ |\   ____\     
-- \|___ \  \_\ \  \|\  \ \  \|\  \     \ \  \___|\ \   __/|\ \  \\ \  \ \   __/|\ \  \|\  \ \  \|\  \|___ \  \_\ \  \ \  \|\  \ \  \\ \  \       \ \  \_|\ \ \   __/|\ \  \___|_        \ \  \___|\ \  \|\  \ \  \\\  \ \  \___|_  ____________\ \  \___|\ \  \    \ \   __/|\ \  \___|_    
--      \ \  \ \ \  \\\  \ \   ____\     \ \  \  __\ \  \_|/_\ \  \\ \  \ \  \_|/_\ \   _  _\ \   __  \   \ \  \ \ \  \ \  \\\  \ \  \\ \  \       \ \  \ \\ \ \  \_|/_\ \_____  \        \ \_____  \ \  \\\  \ \  \\\  \ \_____  \|\____________\ \  \    \ \  \    \ \  \_|/_\ \_____  \   
--       \ \  \ \ \  \\\  \ \  \___|      \ \  \|\  \ \  \_|\ \ \  \\ \  \ \  \_|\ \ \  \\  \\ \  \ \  \   \ \  \ \ \  \ \  \\\  \ \  \\ \  \       \ \  \_\\ \ \  \_|\ \|____|\  \        \|____|\  \ \  \\\  \ \  \\\  \|____|\  \|____________|\ \  \____\ \  \____\ \  \_|\ \|____|\  \  
--        \ \__\ \ \_______\ \__\          \ \_______\ \_______\ \__\\ \__\ \_______\ \__\\ _\\ \__\ \__\   \ \__\ \ \__\ \_______\ \__\\ \__\       \ \_______\ \_______\____\_\  \         ____\_\  \ \_______\ \_______\____\_\  \              \ \_______\ \_______\ \_______\____\_\  \ 
--         \|__|  \|_______|\|__|           \|_______|\|_______|\|__| \|__|\|_______|\|__|\|__|\|__|\|__|    \|__|  \|__|\|_______|\|__| \|__|        \|_______|\|_______|\_________\       |\_________\|_______|\|_______|\_________\              \|_______|\|_______|\|_______|\_________\
--                                                                                                                                                                        \|_________|       \|_________|                  \|_________|                                           \|_________|																																																											  


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.my_package_2.all; 
use work.my_package.all; 


entity aes_top is
    Port (
        clk     : in std_logic;
	rstn    : in std_logic;
        key_in  : in std_logic_vector(127 downto 0);
        key_out : out std_logic_vector(127 downto 0);
	key_select : in integer
    );
end aes_top;

architecture Behavioral of aes_top is
    signal sbox_data	: std_logic_vector(31 downto 0);
    signal sbox_address	: std_logic_vector(31 downto 0);

begin
    key_expansion_inst : entity work.Key_Expansion
    port map (
		clk 	=> clk,
		rstn 	=> rstn,
        key_in  => key_in,
        w0_sub  => sbox_data,
        adress  => sbox_address,
        key_out => key_out,
	    key_select => key_select,
		Gen_key => open
    );

    -- Instanciation de 4 ROM SBOX
    SBOX: for i in 0 to 3 generate
        SBOX_i: entity work.rom_sbox
        port map (
            clk     => clk,
            address => sbox_address(i*8+7 downto i*8),
            data    => sbox_data(i*8+7 downto i*8)
        );
    end generate;

end Behavioral;

