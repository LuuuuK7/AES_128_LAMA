-----------------------------------------------------
-- testbench dechiffrement
-----------------------------------------------------
-- Auteur : Groupe LAMA
-- Date   : fevrier 2023
------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
use work.package_dechiffrement;


entity tb_dechiffrement is
end tb_dechiffrement;

architecture testbench of tb_dechiffrement is
  --Test InvShiftRow
  variable a : array_state;
  a(0,0) <= 

end;